module FILENAME (
  
);
  

endmodule
